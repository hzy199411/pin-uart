/*

Copyright (c) 2023 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`resetall
`timescale 1ns / 1ps
`default_nettype none

/*
 * 
 */
module fpga
(
output wire A4,
output wire A5,
output wire A6,
output wire A7,
output wire A21,
output wire A22,
output wire A24,
output wire A25,
output wire AA1,
output wire AA2,
output wire AA4,
output wire AA5,
output wire AA6,
output wire AA7,
output wire AA9,
output wire AA10,
output wire AA11,
output wire AA12,
output wire AB2,
output wire AB3,
output wire AB4,
output wire AB5,
output wire AB7,
output wire AB8,
output wire AB9,
output wire AB10,
output wire AB12,
output wire AB13,
output wire AC1,
output wire AC2,
output wire AC3,
output wire AC5,
output wire AC6,
output wire AC7,
output wire AC8,
output wire AC10,
output wire AC11,
output wire AC12,
output wire AC13,
output wire AD1,
output wire AD4,
output wire AD5,
output wire AD6,
output wire AD8,
output wire AD9,
output wire AD10,
output wire AD11,
output wire AE1,
output wire AE2,
output wire AE3,
output wire AE4,
output wire AE6,
output wire AE7,
output wire AE8,
output wire AE9,
output wire AE11,
output wire AE12,
output wire AF1,
output wire AF2,
output wire AF4,
output wire AF5,
output wire AF6,
output wire AF7,
output wire AF9,
output wire AF10,
output wire AF11,
output wire AF12,
output wire AG2,
output wire AG3,
output wire AG4,
output wire AG5,
output wire AG7,
output wire AG8,
output wire AG9,
output wire AG10,
output wire AG12,
output wire AG13,
output wire AH1,
output wire AH2,
output wire AH5,
output wire AH6,
output wire AH7,
output wire AH8,
output wire AH10,
output wire AH11,
output wire AH12,
output wire AH13,
output wire AH18,
output wire AH24,
output wire AJ1,
output wire AJ3,
output wire AJ4,
output wire AJ5,
output wire AJ6,
output wire AJ8,
output wire AJ9,
output wire AJ10,
output wire AJ11,
output wire AJ13,
output wire AJ18,
output wire AJ19,
output wire AJ23,
output wire AJ24,
output wire AJ25,
output wire AJ26,
output wire AK1,
output wire AK2,
output wire AK3,
output wire AK4,
output wire AK6,
output wire AK7,
output wire AK8,
output wire AK9,
output wire AK11,
output wire AK12,
output wire AK13,
output wire AK14,
output wire AK17,
output wire AK18,
output wire AK19,
output wire AK21,
output wire AK22,
output wire AK24,
output wire AK27,
output wire AK28,
output wire AK29,
output wire AK30,
output wire AL1,
output wire AL2,
output wire AL4,
output wire AL5,
output wire AL6,
output wire AL7,
output wire AL9,
output wire AL10,
output wire AL11,
output wire AL12,
output wire AL14,
output wire AL17,
output wire AL19,
output wire AL20,
output wire AL21,
output wire AL22,
output wire AL24,
output wire AL25,
output wire AL26,
output wire AL27,
output wire AL29,
output wire AL30,
output wire AM2,
output wire AM3,
output wire AM4,
output wire AM5,
output wire AM7,
output wire AM8,
output wire AM9,
output wire AM10,
output wire AM12,
output wire AM13,
output wire AM17,
output wire AM18,
output wire AM19,
output wire AM20,
output wire AM22,
output wire AM23,
output wire AM24,
output wire AM25,
output wire AM27,
output wire AM29,
output wire AM30,
output wire AN1,
output wire AN2,
output wire AN5,
output wire AN6,
output wire AN7,
output wire AN8,
output wire AN10,
output wire AN11,
output wire AN12,
output wire AN13,
output wire AN17,
output wire AN18,
output wire AN20,
output wire AN21,
output wire AN22,
output wire AN23,
output wire AN25,
output wire AN27,
output wire AN28,
output wire AN30,
output wire AP1,
output wire AP3,
output wire AP4,
output wire AP5,
output wire AP6,
output wire AP8,
output wire AP9,
output wire AP10,
output wire AP11,
output wire AP13,
output wire AP18,
output wire AP19,
output wire AP20,
output wire AP21,
output wire AP23,
output wire AP24,
output wire AP25,
output wire AP26,
output wire AP28,
output wire AP29,
output wire AP30,
output wire AR1,
output wire AR2,
output wire AR3,
output wire AR4,
output wire AR6,
output wire AR7,
output wire AR8,
output wire AR9,
output wire AR11,
output wire AR12,
output wire AR13,
output wire AR16,
output wire AR17,
output wire AR18,
output wire AR19,
output wire AR21,
output wire AR22,
output wire AR23,
output wire AR24,
output wire AR27,
output wire AR28,
output wire AR29,
output wire AR30,
output wire AT1,
output wire AT2,
output wire AT4,
output wire AT5,
output wire AT6,
output wire AT7,
output wire AT9,
output wire AT10,
output wire AT11,
output wire AT12,
output wire AT16,
output wire AT17,
output wire AT19,
output wire AT20,
output wire AT21,
output wire AT22,
output wire AT24,
output wire AT25,
output wire AT26,
output wire AT27,
output wire AT29,
output wire AT30,
output wire AT31,
output wire AU2,
output wire AU3,
output wire AU4,
output wire AU5,
output wire AU7,
output wire AU8,
output wire AU9,
output wire AU10,
output wire AU12,
output wire AU13,
output wire AU17,
output wire AU18,
output wire AU19,
output wire AU20,
output wire AU22,
output wire AU23,
output wire AU24,
output wire AU25,
output wire AU27,
output wire AV1,
output wire AV2,
output wire AV5,
output wire AV6,
output wire AV7,
output wire AV8,
output wire AV10,
output wire AV11,
output wire AV12,
output wire AV16,
output wire AV17,
output wire AV18,
output wire AV20,
output wire AV21,
output wire AV22,
output wire AV23,
output wire AV25,
output wire AV26,
output wire AV27,
output wire AW1,
output wire AW3,
output wire AW4,
output wire AW5,
output wire AW6,
output wire AW8,
output wire AW9,
output wire AW10,
output wire AW11,
output wire AW16,
output wire AW18,
output wire AW19,
output wire AW20,
output wire AW21,
output wire AW23,
output wire AW24,
output wire AW25,
output wire AW26,
output wire AY2,
output wire AY3,
output wire AY4,
output wire AY6,
output wire AY7,
output wire AY16,
output wire AY17,
output wire AY18,
output wire AY19,
output wire AY21,
output wire AY22,
output wire AY23,
output wire AY24,
output wire AY26,
output wire AY27,
output wire B2,
output wire B3,
output wire B4,
output wire B5,
output wire B7,
output wire B22,
output wire B23,
output wire B24,
output wire B25,
output wire BA2,
output wire BA4,
output wire BA5,
output wire BA17,
output wire BA19,
output wire BA20,
output wire BA22,
output wire BA24,
output wire BA25,
output wire BA26,
output wire BA27,
output wire BB4,
output wire BB5,
output wire BB17,
output wire BB18,
output wire BB19,
output wire BB20,
output wire BB22,
output wire BB23,
output wire BB24,
output wire BB25,
output wire BB27,
output wire C2,
output wire C3,
output wire C5,
output wire C6,
output wire C7,
output wire C8,
output wire C10,
output wire C11,
output wire C21,
output wire C22,
output wire C23,
output wire C25,
output wire C26,
output wire C27,
output wire D1,
output wire D3,
output wire D4,
output wire D5,
output wire D6,
output wire D8,
output wire D9,
output wire D10,
output wire D11,
output wire D13,
output wire D14,
output wire D15,
output wire D21,
output wire D23,
output wire D24,
output wire D25,
output wire D26,
output wire D27,
output wire E1,
output wire E2,
output wire E3,
output wire E4,
output wire E6,
output wire E7,
output wire E8,
output wire E9,
output wire E11,
output wire E12,
output wire E13,
output wire E14,
output wire E16,
output wire E21,
output wire E22,
output wire E23,
output wire E24,
output wire E26,
output wire E27,
output wire F1,
output wire F2,
output wire F4,
output wire F5,
output wire F6,
output wire F7,
output wire F9,
output wire F10,
output wire F11,
output wire F12,
output wire F14,
output wire F15,
output wire F16,
output wire F17,
output wire F21,
output wire F22,
output wire F24,
output wire F25,
output wire F26,
output wire F27,
output wire G2,
output wire G3,
output wire G4,
output wire G5,
output wire G7,
output wire G8,
output wire G9,
output wire G10,
output wire G12,
output wire G13,
output wire G14,
output wire G15,
output wire G17,
output wire G22,
output wire G23,
output wire G24,
output wire G25,
output wire G27,
output wire H1,
output wire H2,
output wire H3,
output wire H5,
output wire H6,
output wire H7,
output wire H8,
output wire H10,
output wire H12,
output wire H13,
output wire H15,
output wire H16,
output wire H17,
output wire H21,
output wire H22,
output wire H23,
output wire H25,
output wire H26,
output wire H27,
output wire H28,
output wire H30,
output wire H31,
output wire J1,
output wire J3,
output wire J4,
output wire J6,
output wire J8,
output wire J9,
output wire J10,
output wire J11,
output wire J13,
output wire J15,
output wire J16,
output wire J21,
output wire J23,
output wire J24,
output wire J25,
output wire J28,
output wire J29,
output wire K1,
output wire K2,
output wire K3,
output wire K4,
output wire K6,
output wire K7,
output wire K8,
output wire K9,
output wire K11,
output wire K12,
output wire K13,
output wire K14,
output wire K17,
output wire K22,
output wire K23,
output wire K24,
output wire K26,
output wire K27,
output wire K28,
output wire K29,
output wire K30,
output wire K31,
output wire L1,
output wire L2,
output wire L4,
output wire L5,
output wire L6,
output wire L7,
output wire L9,
output wire L10,
output wire L11,
output wire L12,
output wire L15,
output wire L16,
output wire L17,
output wire L22,
output wire L24,
output wire L25,
output wire L27,
output wire L29,
output wire L30,
output wire M2,
output wire M3,
output wire M4,
output wire M5,
output wire M7,
output wire M8,
output wire M9,
output wire M10,
output wire M12,
output wire M13,
output wire M14,
output wire M15,
output wire M17,
output wire M18,
output wire M22,
output wire M23,
output wire M24,
output wire M25,
output wire M27,
output wire M28,
output wire M29,
output wire M30,
output wire M31,
output wire N1,
output wire N2,
output wire N3,
output wire N5,
output wire N6,
output wire N7,
output wire N8,
output wire N10,
output wire N11,
output wire N12,
output wire N13,
output wire N15,
output wire N16,
output wire N17,
output wire N18,
output wire N23,
output wire N25,
output wire N26,
output wire N27,
output wire N28,
output wire N30,
output wire P1,
output wire P3,
output wire P4,
output wire P6,
output wire P8,
output wire P9,
output wire P10,
output wire P11,
output wire P13,
output wire P15,
output wire P16,
output wire P18,
output wire P23,
output wire P24,
output wire P25,
output wire P26,
output wire P28,
output wire P29,
output wire P30,
output wire P31,
output wire R1,
output wire R2,
output wire R3,
output wire R4,
output wire R6,
output wire R7,
output wire R8,
output wire R9,
output wire R11,
output wire R12,
output wire R13,
output wire R14,
output wire R16,
output wire R17,
output wire R24,
output wire R26,
output wire R27,
output wire T1,
output wire T2,
output wire T4,
output wire T5,
output wire T6,
output wire T7,
output wire T9,
output wire T10,
output wire T11,
output wire T12,
output wire T23,
output wire U2,
output wire U3,
output wire U4,
output wire U5,
output wire U7,
output wire U8,
output wire U9,
output wire U10,
output wire U12,
output wire V1,
output wire V2,
output wire V3,
output wire V5,
output wire V6,
output wire V7,
output wire V8,
output wire V10,
output wire V11,
output wire V12,
output wire W1,
output wire W3,
output wire W4,
output wire W5,
output wire W6,
output wire W8,
output wire W9,
output wire W10,
output wire W11,
output wire Y1,
output wire Y2,
output wire Y4,
output wire Y6,
output wire Y7,
output wire Y8,
output wire Y9,
output wire Y11,
output wire Y12,
output wire Y13
);

wire clk_int;

s10_confclk u0 (
    .clkout (clk_int)
);

localparam CLK_FREQ = 250000000;
localparam BAUD = 115200;
localparam PRESCALE = CLK_FREQ / BAUD;
localparam CL_PRESCALE = $clog2(PRESCALE);


localparam PIN_COUNT = 658;
localparam GROUP_COUNT = 32;
localparam CL_GROUP_COUNT = $clog2(GROUP_COUNT);

reg shift_rst_reg = 1'b0;
reg [CL_GROUP_COUNT-1:0] group_select_reg = 0;
reg [GROUP_COUNT-1:0] shift_reg = 1'b0;

reg [CL_PRESCALE-1:0] prescale_reg = PRESCALE;
reg [5:0] shift_count_reg = 0;

always @(posedge clk_int) begin
    shift_rst_reg <= 1'b0;
    shift_reg <= 0;

    if (prescale_reg) begin
        prescale_reg <= prescale_reg - 1;
    end else begin
        prescale_reg <= PRESCALE;
        if (shift_count_reg) begin
            shift_count_reg <= shift_count_reg - 1;
            shift_reg[group_select_reg] <= 1'b1;
        end else begin
            shift_count_reg <= 6'h3f;
            shift_rst_reg <= 1'b1;
            if (group_select_reg < GROUP_COUNT) begin
                group_select_reg <= group_select_reg + 1;
            end else begin
                group_select_reg <= 0;
            end
        end
    end
end
pin_uart #(.NAME("A4")) pin_A4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[0%GROUP_COUNT]), .out(A4));
pin_uart #(.NAME("A5")) pin_A5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[1%GROUP_COUNT]), .out(A5));
pin_uart #(.NAME("A6")) pin_A6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[2%GROUP_COUNT]), .out(A6));
pin_uart #(.NAME("A7")) pin_A7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[3%GROUP_COUNT]), .out(A7));
pin_uart #(.NAME("A21")) pin_A21_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[4%GROUP_COUNT]), .out(A21));
pin_uart #(.NAME("A22")) pin_A22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[5%GROUP_COUNT]), .out(A22));
pin_uart #(.NAME("A24")) pin_A24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[6%GROUP_COUNT]), .out(A24));
pin_uart #(.NAME("A25")) pin_A25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[7%GROUP_COUNT]), .out(A25));
pin_uart #(.NAME("AA1")) pin_AA1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[8%GROUP_COUNT]), .out(AA1));
pin_uart #(.NAME("AA2")) pin_AA2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[9%GROUP_COUNT]), .out(AA2));
pin_uart #(.NAME("AA4")) pin_AA4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[10%GROUP_COUNT]), .out(AA4));
pin_uart #(.NAME("AA5")) pin_AA5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[11%GROUP_COUNT]), .out(AA5));
pin_uart #(.NAME("AA6")) pin_AA6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[12%GROUP_COUNT]), .out(AA6));
pin_uart #(.NAME("AA7")) pin_AA7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[13%GROUP_COUNT]), .out(AA7));
pin_uart #(.NAME("AA9")) pin_AA9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[14%GROUP_COUNT]), .out(AA9));
pin_uart #(.NAME("AA10")) pin_AA10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[15%GROUP_COUNT]), .out(AA10));
pin_uart #(.NAME("AA11")) pin_AA11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[16%GROUP_COUNT]), .out(AA11));
pin_uart #(.NAME("AA12")) pin_AA12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[17%GROUP_COUNT]), .out(AA12));
pin_uart #(.NAME("AB2")) pin_AB2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[18%GROUP_COUNT]), .out(AB2));
pin_uart #(.NAME("AB3")) pin_AB3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[19%GROUP_COUNT]), .out(AB3));
pin_uart #(.NAME("AB4")) pin_AB4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[20%GROUP_COUNT]), .out(AB4));
pin_uart #(.NAME("AB5")) pin_AB5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[21%GROUP_COUNT]), .out(AB5));
pin_uart #(.NAME("AB7")) pin_AB7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[22%GROUP_COUNT]), .out(AB7));
pin_uart #(.NAME("AB8")) pin_AB8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[23%GROUP_COUNT]), .out(AB8));
pin_uart #(.NAME("AB9")) pin_AB9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[24%GROUP_COUNT]), .out(AB9));
pin_uart #(.NAME("AB10")) pin_AB10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[25%GROUP_COUNT]), .out(AB10));
pin_uart #(.NAME("AB12")) pin_AB12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[26%GROUP_COUNT]), .out(AB12));
pin_uart #(.NAME("AB13")) pin_AB13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[27%GROUP_COUNT]), .out(AB13));
pin_uart #(.NAME("AC1")) pin_AC1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[28%GROUP_COUNT]), .out(AC1));
pin_uart #(.NAME("AC2")) pin_AC2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[29%GROUP_COUNT]), .out(AC2));
pin_uart #(.NAME("AC3")) pin_AC3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[30%GROUP_COUNT]), .out(AC3));
pin_uart #(.NAME("AC5")) pin_AC5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[31%GROUP_COUNT]), .out(AC5));
pin_uart #(.NAME("AC6")) pin_AC6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[32%GROUP_COUNT]), .out(AC6));
pin_uart #(.NAME("AC7")) pin_AC7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[33%GROUP_COUNT]), .out(AC7));
pin_uart #(.NAME("AC8")) pin_AC8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[34%GROUP_COUNT]), .out(AC8));
pin_uart #(.NAME("AC10")) pin_AC10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[35%GROUP_COUNT]), .out(AC10));
pin_uart #(.NAME("AC11")) pin_AC11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[36%GROUP_COUNT]), .out(AC11));
pin_uart #(.NAME("AC12")) pin_AC12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[37%GROUP_COUNT]), .out(AC12));
pin_uart #(.NAME("AC13")) pin_AC13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[38%GROUP_COUNT]), .out(AC13));
pin_uart #(.NAME("AD1")) pin_AD1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[39%GROUP_COUNT]), .out(AD1));
pin_uart #(.NAME("AD4")) pin_AD4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[40%GROUP_COUNT]), .out(AD4));
pin_uart #(.NAME("AD5")) pin_AD5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[41%GROUP_COUNT]), .out(AD5));
pin_uart #(.NAME("AD6")) pin_AD6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[42%GROUP_COUNT]), .out(AD6));
pin_uart #(.NAME("AD8")) pin_AD8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[43%GROUP_COUNT]), .out(AD8));
pin_uart #(.NAME("AD9")) pin_AD9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[44%GROUP_COUNT]), .out(AD9));
pin_uart #(.NAME("AD10")) pin_AD10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[45%GROUP_COUNT]), .out(AD10));
pin_uart #(.NAME("AD11")) pin_AD11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[46%GROUP_COUNT]), .out(AD11));
pin_uart #(.NAME("AE1")) pin_AE1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[47%GROUP_COUNT]), .out(AE1));
pin_uart #(.NAME("AE2")) pin_AE2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[48%GROUP_COUNT]), .out(AE2));
pin_uart #(.NAME("AE3")) pin_AE3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[49%GROUP_COUNT]), .out(AE3));
pin_uart #(.NAME("AE4")) pin_AE4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[50%GROUP_COUNT]), .out(AE4));
pin_uart #(.NAME("AE6")) pin_AE6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[51%GROUP_COUNT]), .out(AE6));
pin_uart #(.NAME("AE7")) pin_AE7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[52%GROUP_COUNT]), .out(AE7));
pin_uart #(.NAME("AE8")) pin_AE8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[53%GROUP_COUNT]), .out(AE8));
pin_uart #(.NAME("AE9")) pin_AE9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[54%GROUP_COUNT]), .out(AE9));
pin_uart #(.NAME("AE11")) pin_AE11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[55%GROUP_COUNT]), .out(AE11));
pin_uart #(.NAME("AE12")) pin_AE12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[56%GROUP_COUNT]), .out(AE12));
pin_uart #(.NAME("AF1")) pin_AF1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[57%GROUP_COUNT]), .out(AF1));
pin_uart #(.NAME("AF2")) pin_AF2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[58%GROUP_COUNT]), .out(AF2));
pin_uart #(.NAME("AF4")) pin_AF4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[59%GROUP_COUNT]), .out(AF4));
pin_uart #(.NAME("AF5")) pin_AF5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[60%GROUP_COUNT]), .out(AF5));
pin_uart #(.NAME("AF6")) pin_AF6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[61%GROUP_COUNT]), .out(AF6));
pin_uart #(.NAME("AF7")) pin_AF7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[62%GROUP_COUNT]), .out(AF7));
pin_uart #(.NAME("AF9")) pin_AF9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[63%GROUP_COUNT]), .out(AF9));
pin_uart #(.NAME("AF10")) pin_AF10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[64%GROUP_COUNT]), .out(AF10));
pin_uart #(.NAME("AF11")) pin_AF11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[65%GROUP_COUNT]), .out(AF11));
pin_uart #(.NAME("AF12")) pin_AF12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[66%GROUP_COUNT]), .out(AF12));
pin_uart #(.NAME("AG2")) pin_AG2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[67%GROUP_COUNT]), .out(AG2));
pin_uart #(.NAME("AG3")) pin_AG3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[68%GROUP_COUNT]), .out(AG3));
pin_uart #(.NAME("AG4")) pin_AG4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[69%GROUP_COUNT]), .out(AG4));
pin_uart #(.NAME("AG5")) pin_AG5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[70%GROUP_COUNT]), .out(AG5));
pin_uart #(.NAME("AG7")) pin_AG7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[71%GROUP_COUNT]), .out(AG7));
pin_uart #(.NAME("AG8")) pin_AG8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[72%GROUP_COUNT]), .out(AG8));
pin_uart #(.NAME("AG9")) pin_AG9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[73%GROUP_COUNT]), .out(AG9));
pin_uart #(.NAME("AG10")) pin_AG10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[74%GROUP_COUNT]), .out(AG10));
pin_uart #(.NAME("AG12")) pin_AG12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[75%GROUP_COUNT]), .out(AG12));
pin_uart #(.NAME("AG13")) pin_AG13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[76%GROUP_COUNT]), .out(AG13));
pin_uart #(.NAME("AH1")) pin_AH1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[77%GROUP_COUNT]), .out(AH1));
pin_uart #(.NAME("AH2")) pin_AH2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[78%GROUP_COUNT]), .out(AH2));
pin_uart #(.NAME("AH5")) pin_AH5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[79%GROUP_COUNT]), .out(AH5));
pin_uart #(.NAME("AH6")) pin_AH6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[80%GROUP_COUNT]), .out(AH6));
pin_uart #(.NAME("AH7")) pin_AH7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[81%GROUP_COUNT]), .out(AH7));
pin_uart #(.NAME("AH8")) pin_AH8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[82%GROUP_COUNT]), .out(AH8));
pin_uart #(.NAME("AH10")) pin_AH10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[83%GROUP_COUNT]), .out(AH10));
pin_uart #(.NAME("AH11")) pin_AH11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[84%GROUP_COUNT]), .out(AH11));
pin_uart #(.NAME("AH12")) pin_AH12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[85%GROUP_COUNT]), .out(AH12));
pin_uart #(.NAME("AH13")) pin_AH13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[86%GROUP_COUNT]), .out(AH13));
pin_uart #(.NAME("AH18")) pin_AH18_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[87%GROUP_COUNT]), .out(AH18));
pin_uart #(.NAME("AH24")) pin_AH24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[88%GROUP_COUNT]), .out(AH24));
pin_uart #(.NAME("AJ1")) pin_AJ1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[89%GROUP_COUNT]), .out(AJ1));
pin_uart #(.NAME("AJ3")) pin_AJ3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[90%GROUP_COUNT]), .out(AJ3));
pin_uart #(.NAME("AJ4")) pin_AJ4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[91%GROUP_COUNT]), .out(AJ4));
pin_uart #(.NAME("AJ5")) pin_AJ5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[92%GROUP_COUNT]), .out(AJ5));
pin_uart #(.NAME("AJ6")) pin_AJ6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[93%GROUP_COUNT]), .out(AJ6));
pin_uart #(.NAME("AJ8")) pin_AJ8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[94%GROUP_COUNT]), .out(AJ8));
pin_uart #(.NAME("AJ9")) pin_AJ9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[95%GROUP_COUNT]), .out(AJ9));
pin_uart #(.NAME("AJ10")) pin_AJ10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[96%GROUP_COUNT]), .out(AJ10));
pin_uart #(.NAME("AJ11")) pin_AJ11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[97%GROUP_COUNT]), .out(AJ11));
pin_uart #(.NAME("AJ13")) pin_AJ13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[98%GROUP_COUNT]), .out(AJ13));
pin_uart #(.NAME("AJ18")) pin_AJ18_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[99%GROUP_COUNT]), .out(AJ18));
pin_uart #(.NAME("AJ19")) pin_AJ19_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[100%GROUP_COUNT]), .out(AJ19));
pin_uart #(.NAME("AJ23")) pin_AJ23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[101%GROUP_COUNT]), .out(AJ23));
pin_uart #(.NAME("AJ24")) pin_AJ24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[102%GROUP_COUNT]), .out(AJ24));
pin_uart #(.NAME("AJ25")) pin_AJ25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[103%GROUP_COUNT]), .out(AJ25));
pin_uart #(.NAME("AJ26")) pin_AJ26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[104%GROUP_COUNT]), .out(AJ26));
pin_uart #(.NAME("AK1")) pin_AK1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[105%GROUP_COUNT]), .out(AK1));
pin_uart #(.NAME("AK2")) pin_AK2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[106%GROUP_COUNT]), .out(AK2));
pin_uart #(.NAME("AK3")) pin_AK3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[107%GROUP_COUNT]), .out(AK3));
pin_uart #(.NAME("AK4")) pin_AK4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[108%GROUP_COUNT]), .out(AK4));
pin_uart #(.NAME("AK6")) pin_AK6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[109%GROUP_COUNT]), .out(AK6));
pin_uart #(.NAME("AK7")) pin_AK7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[110%GROUP_COUNT]), .out(AK7));
pin_uart #(.NAME("AK8")) pin_AK8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[111%GROUP_COUNT]), .out(AK8));
pin_uart #(.NAME("AK9")) pin_AK9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[112%GROUP_COUNT]), .out(AK9));
pin_uart #(.NAME("AK11")) pin_AK11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[113%GROUP_COUNT]), .out(AK11));
pin_uart #(.NAME("AK12")) pin_AK12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[114%GROUP_COUNT]), .out(AK12));
pin_uart #(.NAME("AK13")) pin_AK13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[115%GROUP_COUNT]), .out(AK13));
pin_uart #(.NAME("AK14")) pin_AK14_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[116%GROUP_COUNT]), .out(AK14));
pin_uart #(.NAME("AK17")) pin_AK17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[117%GROUP_COUNT]), .out(AK17));
pin_uart #(.NAME("AK18")) pin_AK18_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[118%GROUP_COUNT]), .out(AK18));
pin_uart #(.NAME("AK19")) pin_AK19_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[119%GROUP_COUNT]), .out(AK19));
pin_uart #(.NAME("AK21")) pin_AK21_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[120%GROUP_COUNT]), .out(AK21));
pin_uart #(.NAME("AK22")) pin_AK22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[121%GROUP_COUNT]), .out(AK22));
pin_uart #(.NAME("AK24")) pin_AK24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[122%GROUP_COUNT]), .out(AK24));
pin_uart #(.NAME("AK27")) pin_AK27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[123%GROUP_COUNT]), .out(AK27));
pin_uart #(.NAME("AK28")) pin_AK28_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[124%GROUP_COUNT]), .out(AK28));
pin_uart #(.NAME("AK29")) pin_AK29_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[125%GROUP_COUNT]), .out(AK29));
pin_uart #(.NAME("AK30")) pin_AK30_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[126%GROUP_COUNT]), .out(AK30));
pin_uart #(.NAME("AL1")) pin_AL1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[127%GROUP_COUNT]), .out(AL1));
pin_uart #(.NAME("AL2")) pin_AL2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[128%GROUP_COUNT]), .out(AL2));
pin_uart #(.NAME("AL4")) pin_AL4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[129%GROUP_COUNT]), .out(AL4));
pin_uart #(.NAME("AL5")) pin_AL5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[130%GROUP_COUNT]), .out(AL5));
pin_uart #(.NAME("AL6")) pin_AL6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[131%GROUP_COUNT]), .out(AL6));
pin_uart #(.NAME("AL7")) pin_AL7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[132%GROUP_COUNT]), .out(AL7));
pin_uart #(.NAME("AL9")) pin_AL9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[133%GROUP_COUNT]), .out(AL9));
pin_uart #(.NAME("AL10")) pin_AL10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[134%GROUP_COUNT]), .out(AL10));
pin_uart #(.NAME("AL11")) pin_AL11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[135%GROUP_COUNT]), .out(AL11));
pin_uart #(.NAME("AL12")) pin_AL12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[136%GROUP_COUNT]), .out(AL12));
pin_uart #(.NAME("AL14")) pin_AL14_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[137%GROUP_COUNT]), .out(AL14));
pin_uart #(.NAME("AL17")) pin_AL17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[138%GROUP_COUNT]), .out(AL17));
pin_uart #(.NAME("AL19")) pin_AL19_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[139%GROUP_COUNT]), .out(AL19));
pin_uart #(.NAME("AL20")) pin_AL20_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[140%GROUP_COUNT]), .out(AL20));
pin_uart #(.NAME("AL21")) pin_AL21_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[141%GROUP_COUNT]), .out(AL21));
pin_uart #(.NAME("AL22")) pin_AL22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[142%GROUP_COUNT]), .out(AL22));
pin_uart #(.NAME("AL24")) pin_AL24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[143%GROUP_COUNT]), .out(AL24));
pin_uart #(.NAME("AL25")) pin_AL25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[144%GROUP_COUNT]), .out(AL25));
pin_uart #(.NAME("AL26")) pin_AL26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[145%GROUP_COUNT]), .out(AL26));
pin_uart #(.NAME("AL27")) pin_AL27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[146%GROUP_COUNT]), .out(AL27));
pin_uart #(.NAME("AL29")) pin_AL29_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[147%GROUP_COUNT]), .out(AL29));
pin_uart #(.NAME("AL30")) pin_AL30_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[148%GROUP_COUNT]), .out(AL30));
pin_uart #(.NAME("AM2")) pin_AM2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[149%GROUP_COUNT]), .out(AM2));
pin_uart #(.NAME("AM3")) pin_AM3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[150%GROUP_COUNT]), .out(AM3));
pin_uart #(.NAME("AM4")) pin_AM4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[151%GROUP_COUNT]), .out(AM4));
pin_uart #(.NAME("AM5")) pin_AM5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[152%GROUP_COUNT]), .out(AM5));
pin_uart #(.NAME("AM7")) pin_AM7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[153%GROUP_COUNT]), .out(AM7));
pin_uart #(.NAME("AM8")) pin_AM8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[154%GROUP_COUNT]), .out(AM8));
pin_uart #(.NAME("AM9")) pin_AM9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[155%GROUP_COUNT]), .out(AM9));
pin_uart #(.NAME("AM10")) pin_AM10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[156%GROUP_COUNT]), .out(AM10));
pin_uart #(.NAME("AM12")) pin_AM12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[157%GROUP_COUNT]), .out(AM12));
pin_uart #(.NAME("AM13")) pin_AM13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[158%GROUP_COUNT]), .out(AM13));
pin_uart #(.NAME("AM17")) pin_AM17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[159%GROUP_COUNT]), .out(AM17));
pin_uart #(.NAME("AM18")) pin_AM18_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[160%GROUP_COUNT]), .out(AM18));
pin_uart #(.NAME("AM19")) pin_AM19_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[161%GROUP_COUNT]), .out(AM19));
pin_uart #(.NAME("AM20")) pin_AM20_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[162%GROUP_COUNT]), .out(AM20));
pin_uart #(.NAME("AM22")) pin_AM22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[163%GROUP_COUNT]), .out(AM22));
pin_uart #(.NAME("AM23")) pin_AM23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[164%GROUP_COUNT]), .out(AM23));
pin_uart #(.NAME("AM24")) pin_AM24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[165%GROUP_COUNT]), .out(AM24));
pin_uart #(.NAME("AM25")) pin_AM25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[166%GROUP_COUNT]), .out(AM25));
pin_uart #(.NAME("AM27")) pin_AM27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[167%GROUP_COUNT]), .out(AM27));
pin_uart #(.NAME("AM29")) pin_AM29_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[168%GROUP_COUNT]), .out(AM29));
pin_uart #(.NAME("AM30")) pin_AM30_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[169%GROUP_COUNT]), .out(AM30));
pin_uart #(.NAME("AN1")) pin_AN1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[170%GROUP_COUNT]), .out(AN1));
pin_uart #(.NAME("AN2")) pin_AN2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[171%GROUP_COUNT]), .out(AN2));
pin_uart #(.NAME("AN5")) pin_AN5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[172%GROUP_COUNT]), .out(AN5));
pin_uart #(.NAME("AN6")) pin_AN6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[173%GROUP_COUNT]), .out(AN6));
pin_uart #(.NAME("AN7")) pin_AN7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[174%GROUP_COUNT]), .out(AN7));
pin_uart #(.NAME("AN8")) pin_AN8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[175%GROUP_COUNT]), .out(AN8));
pin_uart #(.NAME("AN10")) pin_AN10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[176%GROUP_COUNT]), .out(AN10));
pin_uart #(.NAME("AN11")) pin_AN11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[177%GROUP_COUNT]), .out(AN11));
pin_uart #(.NAME("AN12")) pin_AN12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[178%GROUP_COUNT]), .out(AN12));
pin_uart #(.NAME("AN13")) pin_AN13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[179%GROUP_COUNT]), .out(AN13));
pin_uart #(.NAME("AN17")) pin_AN17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[180%GROUP_COUNT]), .out(AN17));
pin_uart #(.NAME("AN18")) pin_AN18_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[181%GROUP_COUNT]), .out(AN18));
pin_uart #(.NAME("AN20")) pin_AN20_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[182%GROUP_COUNT]), .out(AN20));
pin_uart #(.NAME("AN21")) pin_AN21_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[183%GROUP_COUNT]), .out(AN21));
pin_uart #(.NAME("AN22")) pin_AN22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[184%GROUP_COUNT]), .out(AN22));
pin_uart #(.NAME("AN23")) pin_AN23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[185%GROUP_COUNT]), .out(AN23));
pin_uart #(.NAME("AN25")) pin_AN25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[186%GROUP_COUNT]), .out(AN25));
pin_uart #(.NAME("AN27")) pin_AN27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[187%GROUP_COUNT]), .out(AN27));
pin_uart #(.NAME("AN28")) pin_AN28_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[188%GROUP_COUNT]), .out(AN28));
pin_uart #(.NAME("AN30")) pin_AN30_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[189%GROUP_COUNT]), .out(AN30));
pin_uart #(.NAME("AP1")) pin_AP1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[190%GROUP_COUNT]), .out(AP1));
pin_uart #(.NAME("AP3")) pin_AP3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[191%GROUP_COUNT]), .out(AP3));
pin_uart #(.NAME("AP4")) pin_AP4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[192%GROUP_COUNT]), .out(AP4));
pin_uart #(.NAME("AP5")) pin_AP5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[193%GROUP_COUNT]), .out(AP5));
pin_uart #(.NAME("AP6")) pin_AP6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[194%GROUP_COUNT]), .out(AP6));
pin_uart #(.NAME("AP8")) pin_AP8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[195%GROUP_COUNT]), .out(AP8));
pin_uart #(.NAME("AP9")) pin_AP9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[196%GROUP_COUNT]), .out(AP9));
pin_uart #(.NAME("AP10")) pin_AP10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[197%GROUP_COUNT]), .out(AP10));
pin_uart #(.NAME("AP11")) pin_AP11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[198%GROUP_COUNT]), .out(AP11));
pin_uart #(.NAME("AP13")) pin_AP13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[199%GROUP_COUNT]), .out(AP13));
pin_uart #(.NAME("AP18")) pin_AP18_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[200%GROUP_COUNT]), .out(AP18));
pin_uart #(.NAME("AP19")) pin_AP19_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[201%GROUP_COUNT]), .out(AP19));
pin_uart #(.NAME("AP20")) pin_AP20_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[202%GROUP_COUNT]), .out(AP20));
pin_uart #(.NAME("AP21")) pin_AP21_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[203%GROUP_COUNT]), .out(AP21));
pin_uart #(.NAME("AP23")) pin_AP23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[204%GROUP_COUNT]), .out(AP23));
pin_uart #(.NAME("AP24")) pin_AP24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[205%GROUP_COUNT]), .out(AP24));
pin_uart #(.NAME("AP25")) pin_AP25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[206%GROUP_COUNT]), .out(AP25));
pin_uart #(.NAME("AP26")) pin_AP26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[207%GROUP_COUNT]), .out(AP26));
pin_uart #(.NAME("AP28")) pin_AP28_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[208%GROUP_COUNT]), .out(AP28));
pin_uart #(.NAME("AP29")) pin_AP29_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[209%GROUP_COUNT]), .out(AP29));
pin_uart #(.NAME("AP30")) pin_AP30_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[210%GROUP_COUNT]), .out(AP30));
pin_uart #(.NAME("AR1")) pin_AR1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[211%GROUP_COUNT]), .out(AR1));
pin_uart #(.NAME("AR2")) pin_AR2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[212%GROUP_COUNT]), .out(AR2));
pin_uart #(.NAME("AR3")) pin_AR3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[213%GROUP_COUNT]), .out(AR3));
pin_uart #(.NAME("AR4")) pin_AR4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[214%GROUP_COUNT]), .out(AR4));
pin_uart #(.NAME("AR6")) pin_AR6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[215%GROUP_COUNT]), .out(AR6));
pin_uart #(.NAME("AR7")) pin_AR7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[216%GROUP_COUNT]), .out(AR7));
pin_uart #(.NAME("AR8")) pin_AR8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[217%GROUP_COUNT]), .out(AR8));
pin_uart #(.NAME("AR9")) pin_AR9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[218%GROUP_COUNT]), .out(AR9));
pin_uart #(.NAME("AR11")) pin_AR11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[219%GROUP_COUNT]), .out(AR11));
pin_uart #(.NAME("AR12")) pin_AR12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[220%GROUP_COUNT]), .out(AR12));
pin_uart #(.NAME("AR13")) pin_AR13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[221%GROUP_COUNT]), .out(AR13));
pin_uart #(.NAME("AR16")) pin_AR16_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[222%GROUP_COUNT]), .out(AR16));
pin_uart #(.NAME("AR17")) pin_AR17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[223%GROUP_COUNT]), .out(AR17));
pin_uart #(.NAME("AR18")) pin_AR18_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[224%GROUP_COUNT]), .out(AR18));
pin_uart #(.NAME("AR19")) pin_AR19_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[225%GROUP_COUNT]), .out(AR19));
pin_uart #(.NAME("AR21")) pin_AR21_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[226%GROUP_COUNT]), .out(AR21));
pin_uart #(.NAME("AR22")) pin_AR22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[227%GROUP_COUNT]), .out(AR22));
pin_uart #(.NAME("AR23")) pin_AR23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[228%GROUP_COUNT]), .out(AR23));
pin_uart #(.NAME("AR24")) pin_AR24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[229%GROUP_COUNT]), .out(AR24));
pin_uart #(.NAME("AR27")) pin_AR27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[230%GROUP_COUNT]), .out(AR27));
pin_uart #(.NAME("AR28")) pin_AR28_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[231%GROUP_COUNT]), .out(AR28));
pin_uart #(.NAME("AR29")) pin_AR29_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[232%GROUP_COUNT]), .out(AR29));
pin_uart #(.NAME("AR30")) pin_AR30_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[233%GROUP_COUNT]), .out(AR30));
pin_uart #(.NAME("AT1")) pin_AT1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[234%GROUP_COUNT]), .out(AT1));
pin_uart #(.NAME("AT2")) pin_AT2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[235%GROUP_COUNT]), .out(AT2));
pin_uart #(.NAME("AT4")) pin_AT4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[236%GROUP_COUNT]), .out(AT4));
pin_uart #(.NAME("AT5")) pin_AT5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[237%GROUP_COUNT]), .out(AT5));
pin_uart #(.NAME("AT6")) pin_AT6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[238%GROUP_COUNT]), .out(AT6));
pin_uart #(.NAME("AT7")) pin_AT7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[239%GROUP_COUNT]), .out(AT7));
pin_uart #(.NAME("AT9")) pin_AT9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[240%GROUP_COUNT]), .out(AT9));
pin_uart #(.NAME("AT10")) pin_AT10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[241%GROUP_COUNT]), .out(AT10));
pin_uart #(.NAME("AT11")) pin_AT11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[242%GROUP_COUNT]), .out(AT11));
pin_uart #(.NAME("AT12")) pin_AT12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[243%GROUP_COUNT]), .out(AT12));
pin_uart #(.NAME("AT16")) pin_AT16_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[244%GROUP_COUNT]), .out(AT16));
pin_uart #(.NAME("AT17")) pin_AT17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[245%GROUP_COUNT]), .out(AT17));
pin_uart #(.NAME("AT19")) pin_AT19_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[246%GROUP_COUNT]), .out(AT19));
pin_uart #(.NAME("AT20")) pin_AT20_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[247%GROUP_COUNT]), .out(AT20));
pin_uart #(.NAME("AT21")) pin_AT21_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[248%GROUP_COUNT]), .out(AT21));
pin_uart #(.NAME("AT22")) pin_AT22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[249%GROUP_COUNT]), .out(AT22));
pin_uart #(.NAME("AT24")) pin_AT24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[250%GROUP_COUNT]), .out(AT24));
pin_uart #(.NAME("AT25")) pin_AT25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[251%GROUP_COUNT]), .out(AT25));
pin_uart #(.NAME("AT26")) pin_AT26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[252%GROUP_COUNT]), .out(AT26));
pin_uart #(.NAME("AT27")) pin_AT27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[253%GROUP_COUNT]), .out(AT27));
pin_uart #(.NAME("AT29")) pin_AT29_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[254%GROUP_COUNT]), .out(AT29));
pin_uart #(.NAME("AT30")) pin_AT30_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[255%GROUP_COUNT]), .out(AT30));
pin_uart #(.NAME("AT31")) pin_AT31_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[256%GROUP_COUNT]), .out(AT31));
pin_uart #(.NAME("AU2")) pin_AU2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[257%GROUP_COUNT]), .out(AU2));
pin_uart #(.NAME("AU3")) pin_AU3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[258%GROUP_COUNT]), .out(AU3));
pin_uart #(.NAME("AU4")) pin_AU4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[259%GROUP_COUNT]), .out(AU4));
pin_uart #(.NAME("AU5")) pin_AU5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[260%GROUP_COUNT]), .out(AU5));
pin_uart #(.NAME("AU7")) pin_AU7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[261%GROUP_COUNT]), .out(AU7));
pin_uart #(.NAME("AU8")) pin_AU8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[262%GROUP_COUNT]), .out(AU8));
pin_uart #(.NAME("AU9")) pin_AU9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[263%GROUP_COUNT]), .out(AU9));
pin_uart #(.NAME("AU10")) pin_AU10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[264%GROUP_COUNT]), .out(AU10));
pin_uart #(.NAME("AU12")) pin_AU12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[265%GROUP_COUNT]), .out(AU12));
pin_uart #(.NAME("AU13")) pin_AU13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[266%GROUP_COUNT]), .out(AU13));
pin_uart #(.NAME("AU17")) pin_AU17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[267%GROUP_COUNT]), .out(AU17));
pin_uart #(.NAME("AU18")) pin_AU18_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[268%GROUP_COUNT]), .out(AU18));
pin_uart #(.NAME("AU19")) pin_AU19_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[269%GROUP_COUNT]), .out(AU19));
pin_uart #(.NAME("AU20")) pin_AU20_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[270%GROUP_COUNT]), .out(AU20));
pin_uart #(.NAME("AU22")) pin_AU22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[271%GROUP_COUNT]), .out(AU22));
pin_uart #(.NAME("AU23")) pin_AU23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[272%GROUP_COUNT]), .out(AU23));
pin_uart #(.NAME("AU24")) pin_AU24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[273%GROUP_COUNT]), .out(AU24));
pin_uart #(.NAME("AU25")) pin_AU25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[274%GROUP_COUNT]), .out(AU25));
pin_uart #(.NAME("AU27")) pin_AU27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[275%GROUP_COUNT]), .out(AU27));
pin_uart #(.NAME("AV1")) pin_AV1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[276%GROUP_COUNT]), .out(AV1));
pin_uart #(.NAME("AV2")) pin_AV2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[277%GROUP_COUNT]), .out(AV2));
pin_uart #(.NAME("AV5")) pin_AV5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[278%GROUP_COUNT]), .out(AV5));
pin_uart #(.NAME("AV6")) pin_AV6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[279%GROUP_COUNT]), .out(AV6));
pin_uart #(.NAME("AV7")) pin_AV7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[280%GROUP_COUNT]), .out(AV7));
pin_uart #(.NAME("AV8")) pin_AV8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[281%GROUP_COUNT]), .out(AV8));
pin_uart #(.NAME("AV10")) pin_AV10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[282%GROUP_COUNT]), .out(AV10));
pin_uart #(.NAME("AV11")) pin_AV11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[283%GROUP_COUNT]), .out(AV11));
pin_uart #(.NAME("AV12")) pin_AV12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[284%GROUP_COUNT]), .out(AV12));
pin_uart #(.NAME("AV16")) pin_AV16_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[285%GROUP_COUNT]), .out(AV16));
pin_uart #(.NAME("AV17")) pin_AV17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[286%GROUP_COUNT]), .out(AV17));
pin_uart #(.NAME("AV18")) pin_AV18_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[287%GROUP_COUNT]), .out(AV18));
pin_uart #(.NAME("AV20")) pin_AV20_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[288%GROUP_COUNT]), .out(AV20));
pin_uart #(.NAME("AV21")) pin_AV21_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[289%GROUP_COUNT]), .out(AV21));
pin_uart #(.NAME("AV22")) pin_AV22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[290%GROUP_COUNT]), .out(AV22));
pin_uart #(.NAME("AV23")) pin_AV23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[291%GROUP_COUNT]), .out(AV23));
pin_uart #(.NAME("AV25")) pin_AV25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[292%GROUP_COUNT]), .out(AV25));
pin_uart #(.NAME("AV26")) pin_AV26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[293%GROUP_COUNT]), .out(AV26));
pin_uart #(.NAME("AV27")) pin_AV27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[294%GROUP_COUNT]), .out(AV27));
pin_uart #(.NAME("AW1")) pin_AW1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[295%GROUP_COUNT]), .out(AW1));
pin_uart #(.NAME("AW3")) pin_AW3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[296%GROUP_COUNT]), .out(AW3));
pin_uart #(.NAME("AW4")) pin_AW4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[297%GROUP_COUNT]), .out(AW4));
pin_uart #(.NAME("AW5")) pin_AW5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[298%GROUP_COUNT]), .out(AW5));
pin_uart #(.NAME("AW6")) pin_AW6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[299%GROUP_COUNT]), .out(AW6));
pin_uart #(.NAME("AW8")) pin_AW8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[300%GROUP_COUNT]), .out(AW8));
pin_uart #(.NAME("AW9")) pin_AW9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[301%GROUP_COUNT]), .out(AW9));
pin_uart #(.NAME("AW10")) pin_AW10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[302%GROUP_COUNT]), .out(AW10));
pin_uart #(.NAME("AW11")) pin_AW11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[303%GROUP_COUNT]), .out(AW11));
pin_uart #(.NAME("AW16")) pin_AW16_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[304%GROUP_COUNT]), .out(AW16));
pin_uart #(.NAME("AW18")) pin_AW18_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[305%GROUP_COUNT]), .out(AW18));
pin_uart #(.NAME("AW19")) pin_AW19_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[306%GROUP_COUNT]), .out(AW19));
pin_uart #(.NAME("AW20")) pin_AW20_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[307%GROUP_COUNT]), .out(AW20));
pin_uart #(.NAME("AW21")) pin_AW21_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[308%GROUP_COUNT]), .out(AW21));
pin_uart #(.NAME("AW23")) pin_AW23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[309%GROUP_COUNT]), .out(AW23));
pin_uart #(.NAME("AW24")) pin_AW24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[310%GROUP_COUNT]), .out(AW24));
pin_uart #(.NAME("AW25")) pin_AW25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[311%GROUP_COUNT]), .out(AW25));
pin_uart #(.NAME("AW26")) pin_AW26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[312%GROUP_COUNT]), .out(AW26));
pin_uart #(.NAME("AY2")) pin_AY2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[313%GROUP_COUNT]), .out(AY2));
pin_uart #(.NAME("AY3")) pin_AY3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[314%GROUP_COUNT]), .out(AY3));
pin_uart #(.NAME("AY4")) pin_AY4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[315%GROUP_COUNT]), .out(AY4));
pin_uart #(.NAME("AY6")) pin_AY6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[316%GROUP_COUNT]), .out(AY6));
pin_uart #(.NAME("AY7")) pin_AY7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[317%GROUP_COUNT]), .out(AY7));
pin_uart #(.NAME("AY16")) pin_AY16_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[318%GROUP_COUNT]), .out(AY16));
pin_uart #(.NAME("AY17")) pin_AY17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[319%GROUP_COUNT]), .out(AY17));
pin_uart #(.NAME("AY18")) pin_AY18_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[320%GROUP_COUNT]), .out(AY18));
pin_uart #(.NAME("AY19")) pin_AY19_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[321%GROUP_COUNT]), .out(AY19));
pin_uart #(.NAME("AY21")) pin_AY21_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[322%GROUP_COUNT]), .out(AY21));
pin_uart #(.NAME("AY22")) pin_AY22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[323%GROUP_COUNT]), .out(AY22));
pin_uart #(.NAME("AY23")) pin_AY23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[324%GROUP_COUNT]), .out(AY23));
pin_uart #(.NAME("AY24")) pin_AY24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[325%GROUP_COUNT]), .out(AY24));
pin_uart #(.NAME("AY26")) pin_AY26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[326%GROUP_COUNT]), .out(AY26));
pin_uart #(.NAME("AY27")) pin_AY27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[327%GROUP_COUNT]), .out(AY27));
pin_uart #(.NAME("B2")) pin_B2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[328%GROUP_COUNT]), .out(B2));
pin_uart #(.NAME("B3")) pin_B3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[329%GROUP_COUNT]), .out(B3));
pin_uart #(.NAME("B4")) pin_B4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[330%GROUP_COUNT]), .out(B4));
pin_uart #(.NAME("B5")) pin_B5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[331%GROUP_COUNT]), .out(B5));
pin_uart #(.NAME("B7")) pin_B7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[332%GROUP_COUNT]), .out(B7));
pin_uart #(.NAME("B22")) pin_B22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[333%GROUP_COUNT]), .out(B22));
pin_uart #(.NAME("B23")) pin_B23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[334%GROUP_COUNT]), .out(B23));
pin_uart #(.NAME("B24")) pin_B24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[335%GROUP_COUNT]), .out(B24));
pin_uart #(.NAME("B25")) pin_B25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[336%GROUP_COUNT]), .out(B25));
pin_uart #(.NAME("BA2")) pin_BA2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[337%GROUP_COUNT]), .out(BA2));
pin_uart #(.NAME("BA4")) pin_BA4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[338%GROUP_COUNT]), .out(BA4));
pin_uart #(.NAME("BA5")) pin_BA5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[339%GROUP_COUNT]), .out(BA5));
pin_uart #(.NAME("BA17")) pin_BA17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[340%GROUP_COUNT]), .out(BA17));
pin_uart #(.NAME("BA19")) pin_BA19_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[341%GROUP_COUNT]), .out(BA19));
pin_uart #(.NAME("BA20")) pin_BA20_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[342%GROUP_COUNT]), .out(BA20));
pin_uart #(.NAME("BA22")) pin_BA22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[343%GROUP_COUNT]), .out(BA22));
pin_uart #(.NAME("BA24")) pin_BA24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[344%GROUP_COUNT]), .out(BA24));
pin_uart #(.NAME("BA25")) pin_BA25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[345%GROUP_COUNT]), .out(BA25));
pin_uart #(.NAME("BA26")) pin_BA26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[346%GROUP_COUNT]), .out(BA26));
pin_uart #(.NAME("BA27")) pin_BA27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[347%GROUP_COUNT]), .out(BA27));
pin_uart #(.NAME("BB4")) pin_BB4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[348%GROUP_COUNT]), .out(BB4));
pin_uart #(.NAME("BB5")) pin_BB5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[349%GROUP_COUNT]), .out(BB5));
pin_uart #(.NAME("BB17")) pin_BB17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[350%GROUP_COUNT]), .out(BB17));
pin_uart #(.NAME("BB18")) pin_BB18_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[351%GROUP_COUNT]), .out(BB18));
pin_uart #(.NAME("BB19")) pin_BB19_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[352%GROUP_COUNT]), .out(BB19));
pin_uart #(.NAME("BB20")) pin_BB20_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[353%GROUP_COUNT]), .out(BB20));
pin_uart #(.NAME("BB22")) pin_BB22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[354%GROUP_COUNT]), .out(BB22));
pin_uart #(.NAME("BB23")) pin_BB23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[355%GROUP_COUNT]), .out(BB23));
pin_uart #(.NAME("BB24")) pin_BB24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[356%GROUP_COUNT]), .out(BB24));
pin_uart #(.NAME("BB25")) pin_BB25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[357%GROUP_COUNT]), .out(BB25));
pin_uart #(.NAME("BB27")) pin_BB27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[358%GROUP_COUNT]), .out(BB27));
pin_uart #(.NAME("C2")) pin_C2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[359%GROUP_COUNT]), .out(C2));
pin_uart #(.NAME("C3")) pin_C3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[360%GROUP_COUNT]), .out(C3));
pin_uart #(.NAME("C5")) pin_C5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[361%GROUP_COUNT]), .out(C5));
pin_uart #(.NAME("C6")) pin_C6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[362%GROUP_COUNT]), .out(C6));
pin_uart #(.NAME("C7")) pin_C7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[363%GROUP_COUNT]), .out(C7));
pin_uart #(.NAME("C8")) pin_C8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[364%GROUP_COUNT]), .out(C8));
pin_uart #(.NAME("C10")) pin_C10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[365%GROUP_COUNT]), .out(C10));
pin_uart #(.NAME("C11")) pin_C11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[366%GROUP_COUNT]), .out(C11));
pin_uart #(.NAME("C21")) pin_C21_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[367%GROUP_COUNT]), .out(C21));
pin_uart #(.NAME("C22")) pin_C22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[368%GROUP_COUNT]), .out(C22));
pin_uart #(.NAME("C23")) pin_C23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[369%GROUP_COUNT]), .out(C23));
pin_uart #(.NAME("C25")) pin_C25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[370%GROUP_COUNT]), .out(C25));
pin_uart #(.NAME("C26")) pin_C26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[371%GROUP_COUNT]), .out(C26));
pin_uart #(.NAME("C27")) pin_C27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[372%GROUP_COUNT]), .out(C27));
pin_uart #(.NAME("D1")) pin_D1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[373%GROUP_COUNT]), .out(D1));
pin_uart #(.NAME("D3")) pin_D3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[374%GROUP_COUNT]), .out(D3));
pin_uart #(.NAME("D4")) pin_D4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[375%GROUP_COUNT]), .out(D4));
pin_uart #(.NAME("D5")) pin_D5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[376%GROUP_COUNT]), .out(D5));
pin_uart #(.NAME("D6")) pin_D6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[377%GROUP_COUNT]), .out(D6));
pin_uart #(.NAME("D8")) pin_D8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[378%GROUP_COUNT]), .out(D8));
pin_uart #(.NAME("D9")) pin_D9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[379%GROUP_COUNT]), .out(D9));
pin_uart #(.NAME("D10")) pin_D10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[380%GROUP_COUNT]), .out(D10));
pin_uart #(.NAME("D11")) pin_D11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[381%GROUP_COUNT]), .out(D11));
pin_uart #(.NAME("D13")) pin_D13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[382%GROUP_COUNT]), .out(D13));
pin_uart #(.NAME("D14")) pin_D14_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[383%GROUP_COUNT]), .out(D14));
pin_uart #(.NAME("D15")) pin_D15_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[384%GROUP_COUNT]), .out(D15));
pin_uart #(.NAME("D21")) pin_D21_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[385%GROUP_COUNT]), .out(D21));
pin_uart #(.NAME("D23")) pin_D23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[386%GROUP_COUNT]), .out(D23));
pin_uart #(.NAME("D24")) pin_D24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[387%GROUP_COUNT]), .out(D24));
pin_uart #(.NAME("D25")) pin_D25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[388%GROUP_COUNT]), .out(D25));
pin_uart #(.NAME("D26")) pin_D26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[389%GROUP_COUNT]), .out(D26));
pin_uart #(.NAME("D27")) pin_D27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[390%GROUP_COUNT]), .out(D27));
pin_uart #(.NAME("E1")) pin_E1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[391%GROUP_COUNT]), .out(E1));
pin_uart #(.NAME("E2")) pin_E2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[392%GROUP_COUNT]), .out(E2));
pin_uart #(.NAME("E3")) pin_E3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[393%GROUP_COUNT]), .out(E3));
pin_uart #(.NAME("E4")) pin_E4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[394%GROUP_COUNT]), .out(E4));
pin_uart #(.NAME("E6")) pin_E6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[395%GROUP_COUNT]), .out(E6));
pin_uart #(.NAME("E7")) pin_E7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[396%GROUP_COUNT]), .out(E7));
pin_uart #(.NAME("E8")) pin_E8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[397%GROUP_COUNT]), .out(E8));
pin_uart #(.NAME("E9")) pin_E9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[398%GROUP_COUNT]), .out(E9));
pin_uart #(.NAME("E11")) pin_E11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[399%GROUP_COUNT]), .out(E11));
pin_uart #(.NAME("E12")) pin_E12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[400%GROUP_COUNT]), .out(E12));
pin_uart #(.NAME("E13")) pin_E13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[401%GROUP_COUNT]), .out(E13));
pin_uart #(.NAME("E14")) pin_E14_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[402%GROUP_COUNT]), .out(E14));
pin_uart #(.NAME("E16")) pin_E16_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[403%GROUP_COUNT]), .out(E16));
pin_uart #(.NAME("E21")) pin_E21_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[404%GROUP_COUNT]), .out(E21));
pin_uart #(.NAME("E22")) pin_E22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[405%GROUP_COUNT]), .out(E22));
pin_uart #(.NAME("E23")) pin_E23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[406%GROUP_COUNT]), .out(E23));
pin_uart #(.NAME("E24")) pin_E24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[407%GROUP_COUNT]), .out(E24));
pin_uart #(.NAME("E26")) pin_E26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[408%GROUP_COUNT]), .out(E26));
pin_uart #(.NAME("E27")) pin_E27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[409%GROUP_COUNT]), .out(E27));
pin_uart #(.NAME("F1")) pin_F1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[410%GROUP_COUNT]), .out(F1));
pin_uart #(.NAME("F2")) pin_F2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[411%GROUP_COUNT]), .out(F2));
pin_uart #(.NAME("F4")) pin_F4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[412%GROUP_COUNT]), .out(F4));
pin_uart #(.NAME("F5")) pin_F5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[413%GROUP_COUNT]), .out(F5));
pin_uart #(.NAME("F6")) pin_F6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[414%GROUP_COUNT]), .out(F6));
pin_uart #(.NAME("F7")) pin_F7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[415%GROUP_COUNT]), .out(F7));
pin_uart #(.NAME("F9")) pin_F9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[416%GROUP_COUNT]), .out(F9));
pin_uart #(.NAME("F10")) pin_F10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[417%GROUP_COUNT]), .out(F10));
pin_uart #(.NAME("F11")) pin_F11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[418%GROUP_COUNT]), .out(F11));
pin_uart #(.NAME("F12")) pin_F12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[419%GROUP_COUNT]), .out(F12));
pin_uart #(.NAME("F14")) pin_F14_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[420%GROUP_COUNT]), .out(F14));
pin_uart #(.NAME("F15")) pin_F15_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[421%GROUP_COUNT]), .out(F15));
pin_uart #(.NAME("F16")) pin_F16_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[422%GROUP_COUNT]), .out(F16));
pin_uart #(.NAME("F17")) pin_F17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[423%GROUP_COUNT]), .out(F17));
pin_uart #(.NAME("F21")) pin_F21_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[424%GROUP_COUNT]), .out(F21));
pin_uart #(.NAME("F22")) pin_F22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[425%GROUP_COUNT]), .out(F22));
pin_uart #(.NAME("F24")) pin_F24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[426%GROUP_COUNT]), .out(F24));
pin_uart #(.NAME("F25")) pin_F25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[427%GROUP_COUNT]), .out(F25));
pin_uart #(.NAME("F26")) pin_F26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[428%GROUP_COUNT]), .out(F26));
pin_uart #(.NAME("F27")) pin_F27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[429%GROUP_COUNT]), .out(F27));
pin_uart #(.NAME("G2")) pin_G2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[430%GROUP_COUNT]), .out(G2));
pin_uart #(.NAME("G3")) pin_G3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[431%GROUP_COUNT]), .out(G3));
pin_uart #(.NAME("G4")) pin_G4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[432%GROUP_COUNT]), .out(G4));
pin_uart #(.NAME("G5")) pin_G5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[433%GROUP_COUNT]), .out(G5));
pin_uart #(.NAME("G7")) pin_G7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[434%GROUP_COUNT]), .out(G7));
pin_uart #(.NAME("G8")) pin_G8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[435%GROUP_COUNT]), .out(G8));
pin_uart #(.NAME("G9")) pin_G9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[436%GROUP_COUNT]), .out(G9));
pin_uart #(.NAME("G10")) pin_G10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[437%GROUP_COUNT]), .out(G10));
pin_uart #(.NAME("G12")) pin_G12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[438%GROUP_COUNT]), .out(G12));
pin_uart #(.NAME("G13")) pin_G13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[439%GROUP_COUNT]), .out(G13));
pin_uart #(.NAME("G14")) pin_G14_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[440%GROUP_COUNT]), .out(G14));
pin_uart #(.NAME("G15")) pin_G15_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[441%GROUP_COUNT]), .out(G15));
pin_uart #(.NAME("G17")) pin_G17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[442%GROUP_COUNT]), .out(G17));
pin_uart #(.NAME("G22")) pin_G22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[443%GROUP_COUNT]), .out(G22));
pin_uart #(.NAME("G23")) pin_G23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[444%GROUP_COUNT]), .out(G23));
pin_uart #(.NAME("G24")) pin_G24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[445%GROUP_COUNT]), .out(G24));
pin_uart #(.NAME("G25")) pin_G25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[446%GROUP_COUNT]), .out(G25));
pin_uart #(.NAME("G27")) pin_G27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[447%GROUP_COUNT]), .out(G27));
pin_uart #(.NAME("H1")) pin_H1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[448%GROUP_COUNT]), .out(H1));
pin_uart #(.NAME("H2")) pin_H2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[449%GROUP_COUNT]), .out(H2));
pin_uart #(.NAME("H3")) pin_H3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[450%GROUP_COUNT]), .out(H3));
pin_uart #(.NAME("H5")) pin_H5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[451%GROUP_COUNT]), .out(H5));
pin_uart #(.NAME("H6")) pin_H6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[452%GROUP_COUNT]), .out(H6));
pin_uart #(.NAME("H7")) pin_H7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[453%GROUP_COUNT]), .out(H7));
pin_uart #(.NAME("H8")) pin_H8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[454%GROUP_COUNT]), .out(H8));
pin_uart #(.NAME("H10")) pin_H10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[455%GROUP_COUNT]), .out(H10));
pin_uart #(.NAME("H12")) pin_H12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[456%GROUP_COUNT]), .out(H12));
pin_uart #(.NAME("H13")) pin_H13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[457%GROUP_COUNT]), .out(H13));
pin_uart #(.NAME("H15")) pin_H15_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[458%GROUP_COUNT]), .out(H15));
pin_uart #(.NAME("H16")) pin_H16_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[459%GROUP_COUNT]), .out(H16));
pin_uart #(.NAME("H17")) pin_H17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[460%GROUP_COUNT]), .out(H17));
pin_uart #(.NAME("H21")) pin_H21_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[461%GROUP_COUNT]), .out(H21));
pin_uart #(.NAME("H22")) pin_H22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[462%GROUP_COUNT]), .out(H22));
pin_uart #(.NAME("H23")) pin_H23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[463%GROUP_COUNT]), .out(H23));
pin_uart #(.NAME("H25")) pin_H25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[464%GROUP_COUNT]), .out(H25));
pin_uart #(.NAME("H26")) pin_H26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[465%GROUP_COUNT]), .out(H26));
pin_uart #(.NAME("H27")) pin_H27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[466%GROUP_COUNT]), .out(H27));
pin_uart #(.NAME("H28")) pin_H28_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[467%GROUP_COUNT]), .out(H28));
pin_uart #(.NAME("H30")) pin_H30_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[468%GROUP_COUNT]), .out(H30));
pin_uart #(.NAME("H31")) pin_H31_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[469%GROUP_COUNT]), .out(H31));
pin_uart #(.NAME("J1")) pin_J1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[470%GROUP_COUNT]), .out(J1));
pin_uart #(.NAME("J3")) pin_J3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[471%GROUP_COUNT]), .out(J3));
pin_uart #(.NAME("J4")) pin_J4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[472%GROUP_COUNT]), .out(J4));
pin_uart #(.NAME("J6")) pin_J6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[473%GROUP_COUNT]), .out(J6));
pin_uart #(.NAME("J8")) pin_J8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[474%GROUP_COUNT]), .out(J8));
pin_uart #(.NAME("J9")) pin_J9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[475%GROUP_COUNT]), .out(J9));
pin_uart #(.NAME("J10")) pin_J10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[476%GROUP_COUNT]), .out(J10));
pin_uart #(.NAME("J11")) pin_J11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[477%GROUP_COUNT]), .out(J11));
pin_uart #(.NAME("J13")) pin_J13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[478%GROUP_COUNT]), .out(J13));
pin_uart #(.NAME("J15")) pin_J15_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[479%GROUP_COUNT]), .out(J15));
pin_uart #(.NAME("J16")) pin_J16_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[480%GROUP_COUNT]), .out(J16));
pin_uart #(.NAME("J21")) pin_J21_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[481%GROUP_COUNT]), .out(J21));
pin_uart #(.NAME("J23")) pin_J23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[482%GROUP_COUNT]), .out(J23));
pin_uart #(.NAME("J24")) pin_J24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[483%GROUP_COUNT]), .out(J24));
pin_uart #(.NAME("J25")) pin_J25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[484%GROUP_COUNT]), .out(J25));
pin_uart #(.NAME("J28")) pin_J28_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[485%GROUP_COUNT]), .out(J28));
pin_uart #(.NAME("J29")) pin_J29_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[486%GROUP_COUNT]), .out(J29));
pin_uart #(.NAME("K1")) pin_K1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[487%GROUP_COUNT]), .out(K1));
pin_uart #(.NAME("K2")) pin_K2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[488%GROUP_COUNT]), .out(K2));
pin_uart #(.NAME("K3")) pin_K3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[489%GROUP_COUNT]), .out(K3));
pin_uart #(.NAME("K4")) pin_K4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[490%GROUP_COUNT]), .out(K4));
pin_uart #(.NAME("K6")) pin_K6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[491%GROUP_COUNT]), .out(K6));
pin_uart #(.NAME("K7")) pin_K7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[492%GROUP_COUNT]), .out(K7));
pin_uart #(.NAME("K8")) pin_K8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[493%GROUP_COUNT]), .out(K8));
pin_uart #(.NAME("K9")) pin_K9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[494%GROUP_COUNT]), .out(K9));
pin_uart #(.NAME("K11")) pin_K11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[495%GROUP_COUNT]), .out(K11));
pin_uart #(.NAME("K12")) pin_K12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[496%GROUP_COUNT]), .out(K12));
pin_uart #(.NAME("K13")) pin_K13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[497%GROUP_COUNT]), .out(K13));
pin_uart #(.NAME("K14")) pin_K14_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[498%GROUP_COUNT]), .out(K14));
pin_uart #(.NAME("K17")) pin_K17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[499%GROUP_COUNT]), .out(K17));
pin_uart #(.NAME("K22")) pin_K22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[500%GROUP_COUNT]), .out(K22));
pin_uart #(.NAME("K23")) pin_K23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[501%GROUP_COUNT]), .out(K23));
pin_uart #(.NAME("K24")) pin_K24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[502%GROUP_COUNT]), .out(K24));
pin_uart #(.NAME("K26")) pin_K26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[503%GROUP_COUNT]), .out(K26));
pin_uart #(.NAME("K27")) pin_K27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[504%GROUP_COUNT]), .out(K27));
pin_uart #(.NAME("K28")) pin_K28_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[505%GROUP_COUNT]), .out(K28));
pin_uart #(.NAME("K29")) pin_K29_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[506%GROUP_COUNT]), .out(K29));
pin_uart #(.NAME("K30")) pin_K30_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[507%GROUP_COUNT]), .out(K30));
pin_uart #(.NAME("K31")) pin_K31_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[508%GROUP_COUNT]), .out(K31));
pin_uart #(.NAME("L1")) pin_L1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[509%GROUP_COUNT]), .out(L1));
pin_uart #(.NAME("L2")) pin_L2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[510%GROUP_COUNT]), .out(L2));
pin_uart #(.NAME("L4")) pin_L4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[511%GROUP_COUNT]), .out(L4));
pin_uart #(.NAME("L5")) pin_L5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[512%GROUP_COUNT]), .out(L5));
pin_uart #(.NAME("L6")) pin_L6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[513%GROUP_COUNT]), .out(L6));
pin_uart #(.NAME("L7")) pin_L7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[514%GROUP_COUNT]), .out(L7));
pin_uart #(.NAME("L9")) pin_L9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[515%GROUP_COUNT]), .out(L9));
pin_uart #(.NAME("L10")) pin_L10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[516%GROUP_COUNT]), .out(L10));
pin_uart #(.NAME("L11")) pin_L11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[517%GROUP_COUNT]), .out(L11));
pin_uart #(.NAME("L12")) pin_L12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[518%GROUP_COUNT]), .out(L12));
pin_uart #(.NAME("L15")) pin_L15_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[519%GROUP_COUNT]), .out(L15));
pin_uart #(.NAME("L16")) pin_L16_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[520%GROUP_COUNT]), .out(L16));
pin_uart #(.NAME("L17")) pin_L17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[521%GROUP_COUNT]), .out(L17));
pin_uart #(.NAME("L22")) pin_L22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[522%GROUP_COUNT]), .out(L22));
pin_uart #(.NAME("L24")) pin_L24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[523%GROUP_COUNT]), .out(L24));
pin_uart #(.NAME("L25")) pin_L25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[524%GROUP_COUNT]), .out(L25));
pin_uart #(.NAME("L27")) pin_L27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[525%GROUP_COUNT]), .out(L27));
pin_uart #(.NAME("L29")) pin_L29_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[526%GROUP_COUNT]), .out(L29));
pin_uart #(.NAME("L30")) pin_L30_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[527%GROUP_COUNT]), .out(L30));
pin_uart #(.NAME("M2")) pin_M2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[528%GROUP_COUNT]), .out(M2));
pin_uart #(.NAME("M3")) pin_M3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[529%GROUP_COUNT]), .out(M3));
pin_uart #(.NAME("M4")) pin_M4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[530%GROUP_COUNT]), .out(M4));
pin_uart #(.NAME("M5")) pin_M5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[531%GROUP_COUNT]), .out(M5));
pin_uart #(.NAME("M7")) pin_M7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[532%GROUP_COUNT]), .out(M7));
pin_uart #(.NAME("M8")) pin_M8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[533%GROUP_COUNT]), .out(M8));
pin_uart #(.NAME("M9")) pin_M9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[534%GROUP_COUNT]), .out(M9));
pin_uart #(.NAME("M10")) pin_M10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[535%GROUP_COUNT]), .out(M10));
pin_uart #(.NAME("M12")) pin_M12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[536%GROUP_COUNT]), .out(M12));
pin_uart #(.NAME("M13")) pin_M13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[537%GROUP_COUNT]), .out(M13));
pin_uart #(.NAME("M14")) pin_M14_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[538%GROUP_COUNT]), .out(M14));
pin_uart #(.NAME("M15")) pin_M15_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[539%GROUP_COUNT]), .out(M15));
pin_uart #(.NAME("M17")) pin_M17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[540%GROUP_COUNT]), .out(M17));
pin_uart #(.NAME("M18")) pin_M18_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[541%GROUP_COUNT]), .out(M18));
pin_uart #(.NAME("M22")) pin_M22_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[542%GROUP_COUNT]), .out(M22));
pin_uart #(.NAME("M23")) pin_M23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[543%GROUP_COUNT]), .out(M23));
pin_uart #(.NAME("M24")) pin_M24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[544%GROUP_COUNT]), .out(M24));
pin_uart #(.NAME("M25")) pin_M25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[545%GROUP_COUNT]), .out(M25));
pin_uart #(.NAME("M27")) pin_M27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[546%GROUP_COUNT]), .out(M27));
pin_uart #(.NAME("M28")) pin_M28_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[547%GROUP_COUNT]), .out(M28));
pin_uart #(.NAME("M29")) pin_M29_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[548%GROUP_COUNT]), .out(M29));
pin_uart #(.NAME("M30")) pin_M30_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[549%GROUP_COUNT]), .out(M30));
pin_uart #(.NAME("M31")) pin_M31_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[550%GROUP_COUNT]), .out(M31));
pin_uart #(.NAME("N1")) pin_N1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[551%GROUP_COUNT]), .out(N1));
pin_uart #(.NAME("N2")) pin_N2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[552%GROUP_COUNT]), .out(N2));
pin_uart #(.NAME("N3")) pin_N3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[553%GROUP_COUNT]), .out(N3));
pin_uart #(.NAME("N5")) pin_N5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[554%GROUP_COUNT]), .out(N5));
pin_uart #(.NAME("N6")) pin_N6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[555%GROUP_COUNT]), .out(N6));
pin_uart #(.NAME("N7")) pin_N7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[556%GROUP_COUNT]), .out(N7));
pin_uart #(.NAME("N8")) pin_N8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[557%GROUP_COUNT]), .out(N8));
pin_uart #(.NAME("N10")) pin_N10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[558%GROUP_COUNT]), .out(N10));
pin_uart #(.NAME("N11")) pin_N11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[559%GROUP_COUNT]), .out(N11));
pin_uart #(.NAME("N12")) pin_N12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[560%GROUP_COUNT]), .out(N12));
pin_uart #(.NAME("N13")) pin_N13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[561%GROUP_COUNT]), .out(N13));
pin_uart #(.NAME("N15")) pin_N15_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[562%GROUP_COUNT]), .out(N15));
pin_uart #(.NAME("N16")) pin_N16_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[563%GROUP_COUNT]), .out(N16));
pin_uart #(.NAME("N17")) pin_N17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[564%GROUP_COUNT]), .out(N17));
pin_uart #(.NAME("N18")) pin_N18_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[565%GROUP_COUNT]), .out(N18));
pin_uart #(.NAME("N23")) pin_N23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[566%GROUP_COUNT]), .out(N23));
pin_uart #(.NAME("N25")) pin_N25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[567%GROUP_COUNT]), .out(N25));
pin_uart #(.NAME("N26")) pin_N26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[568%GROUP_COUNT]), .out(N26));
pin_uart #(.NAME("N27")) pin_N27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[569%GROUP_COUNT]), .out(N27));
pin_uart #(.NAME("N28")) pin_N28_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[570%GROUP_COUNT]), .out(N28));
pin_uart #(.NAME("N30")) pin_N30_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[571%GROUP_COUNT]), .out(N30));
pin_uart #(.NAME("P1")) pin_P1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[572%GROUP_COUNT]), .out(P1));
pin_uart #(.NAME("P3")) pin_P3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[573%GROUP_COUNT]), .out(P3));
pin_uart #(.NAME("P4")) pin_P4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[574%GROUP_COUNT]), .out(P4));
pin_uart #(.NAME("P6")) pin_P6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[575%GROUP_COUNT]), .out(P6));
pin_uart #(.NAME("P8")) pin_P8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[576%GROUP_COUNT]), .out(P8));
pin_uart #(.NAME("P9")) pin_P9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[577%GROUP_COUNT]), .out(P9));
pin_uart #(.NAME("P10")) pin_P10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[578%GROUP_COUNT]), .out(P10));
pin_uart #(.NAME("P11")) pin_P11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[579%GROUP_COUNT]), .out(P11));
pin_uart #(.NAME("P13")) pin_P13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[580%GROUP_COUNT]), .out(P13));
pin_uart #(.NAME("P15")) pin_P15_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[581%GROUP_COUNT]), .out(P15));
pin_uart #(.NAME("P16")) pin_P16_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[582%GROUP_COUNT]), .out(P16));
pin_uart #(.NAME("P18")) pin_P18_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[583%GROUP_COUNT]), .out(P18));
pin_uart #(.NAME("P23")) pin_P23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[584%GROUP_COUNT]), .out(P23));
pin_uart #(.NAME("P24")) pin_P24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[585%GROUP_COUNT]), .out(P24));
pin_uart #(.NAME("P25")) pin_P25_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[586%GROUP_COUNT]), .out(P25));
pin_uart #(.NAME("P26")) pin_P26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[587%GROUP_COUNT]), .out(P26));
pin_uart #(.NAME("P28")) pin_P28_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[588%GROUP_COUNT]), .out(P28));
pin_uart #(.NAME("P29")) pin_P29_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[589%GROUP_COUNT]), .out(P29));
pin_uart #(.NAME("P30")) pin_P30_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[590%GROUP_COUNT]), .out(P30));
pin_uart #(.NAME("P31")) pin_P31_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[591%GROUP_COUNT]), .out(P31));
pin_uart #(.NAME("R1")) pin_R1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[592%GROUP_COUNT]), .out(R1));
pin_uart #(.NAME("R2")) pin_R2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[593%GROUP_COUNT]), .out(R2));
pin_uart #(.NAME("R3")) pin_R3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[594%GROUP_COUNT]), .out(R3));
pin_uart #(.NAME("R4")) pin_R4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[595%GROUP_COUNT]), .out(R4));
pin_uart #(.NAME("R6")) pin_R6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[596%GROUP_COUNT]), .out(R6));
pin_uart #(.NAME("R7")) pin_R7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[597%GROUP_COUNT]), .out(R7));
pin_uart #(.NAME("R8")) pin_R8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[598%GROUP_COUNT]), .out(R8));
pin_uart #(.NAME("R9")) pin_R9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[599%GROUP_COUNT]), .out(R9));
pin_uart #(.NAME("R11")) pin_R11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[600%GROUP_COUNT]), .out(R11));
pin_uart #(.NAME("R12")) pin_R12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[601%GROUP_COUNT]), .out(R12));
pin_uart #(.NAME("R13")) pin_R13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[602%GROUP_COUNT]), .out(R13));
pin_uart #(.NAME("R14")) pin_R14_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[603%GROUP_COUNT]), .out(R14));
pin_uart #(.NAME("R16")) pin_R16_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[604%GROUP_COUNT]), .out(R16));
pin_uart #(.NAME("R17")) pin_R17_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[605%GROUP_COUNT]), .out(R17));
pin_uart #(.NAME("R24")) pin_R24_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[606%GROUP_COUNT]), .out(R24));
pin_uart #(.NAME("R26")) pin_R26_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[607%GROUP_COUNT]), .out(R26));
pin_uart #(.NAME("R27")) pin_R27_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[608%GROUP_COUNT]), .out(R27));
pin_uart #(.NAME("T1")) pin_T1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[609%GROUP_COUNT]), .out(T1));
pin_uart #(.NAME("T2")) pin_T2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[610%GROUP_COUNT]), .out(T2));
pin_uart #(.NAME("T4")) pin_T4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[611%GROUP_COUNT]), .out(T4));
pin_uart #(.NAME("T5")) pin_T5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[612%GROUP_COUNT]), .out(T5));
pin_uart #(.NAME("T6")) pin_T6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[613%GROUP_COUNT]), .out(T6));
pin_uart #(.NAME("T7")) pin_T7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[614%GROUP_COUNT]), .out(T7));
pin_uart #(.NAME("T9")) pin_T9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[615%GROUP_COUNT]), .out(T9));
pin_uart #(.NAME("T10")) pin_T10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[616%GROUP_COUNT]), .out(T10));
pin_uart #(.NAME("T11")) pin_T11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[617%GROUP_COUNT]), .out(T11));
pin_uart #(.NAME("T12")) pin_T12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[618%GROUP_COUNT]), .out(T12));
pin_uart #(.NAME("T23")) pin_T23_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[619%GROUP_COUNT]), .out(T23));
pin_uart #(.NAME("U2")) pin_U2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[620%GROUP_COUNT]), .out(U2));
pin_uart #(.NAME("U3")) pin_U3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[621%GROUP_COUNT]), .out(U3));
pin_uart #(.NAME("U4")) pin_U4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[622%GROUP_COUNT]), .out(U4));
pin_uart #(.NAME("U5")) pin_U5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[623%GROUP_COUNT]), .out(U5));
pin_uart #(.NAME("U7")) pin_U7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[624%GROUP_COUNT]), .out(U7));
pin_uart #(.NAME("U8")) pin_U8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[625%GROUP_COUNT]), .out(U8));
pin_uart #(.NAME("U9")) pin_U9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[626%GROUP_COUNT]), .out(U9));
pin_uart #(.NAME("U10")) pin_U10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[627%GROUP_COUNT]), .out(U10));
pin_uart #(.NAME("U12")) pin_U12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[628%GROUP_COUNT]), .out(U12));
pin_uart #(.NAME("V1")) pin_V1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[629%GROUP_COUNT]), .out(V1));
pin_uart #(.NAME("V2")) pin_V2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[630%GROUP_COUNT]), .out(V2));
pin_uart #(.NAME("V3")) pin_V3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[631%GROUP_COUNT]), .out(V3));
pin_uart #(.NAME("V5")) pin_V5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[632%GROUP_COUNT]), .out(V5));
pin_uart #(.NAME("V6")) pin_V6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[633%GROUP_COUNT]), .out(V6));
pin_uart #(.NAME("V7")) pin_V7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[634%GROUP_COUNT]), .out(V7));
pin_uart #(.NAME("V8")) pin_V8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[635%GROUP_COUNT]), .out(V8));
pin_uart #(.NAME("V10")) pin_V10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[636%GROUP_COUNT]), .out(V10));
pin_uart #(.NAME("V11")) pin_V11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[637%GROUP_COUNT]), .out(V11));
pin_uart #(.NAME("V12")) pin_V12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[638%GROUP_COUNT]), .out(V12));
pin_uart #(.NAME("W1")) pin_W1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[639%GROUP_COUNT]), .out(W1));
pin_uart #(.NAME("W3")) pin_W3_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[640%GROUP_COUNT]), .out(W3));
pin_uart #(.NAME("W4")) pin_W4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[641%GROUP_COUNT]), .out(W4));
pin_uart #(.NAME("W5")) pin_W5_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[642%GROUP_COUNT]), .out(W5));
pin_uart #(.NAME("W6")) pin_W6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[643%GROUP_COUNT]), .out(W6));
pin_uart #(.NAME("W8")) pin_W8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[644%GROUP_COUNT]), .out(W8));
pin_uart #(.NAME("W9")) pin_W9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[645%GROUP_COUNT]), .out(W9));
pin_uart #(.NAME("W10")) pin_W10_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[646%GROUP_COUNT]), .out(W10));
pin_uart #(.NAME("W11")) pin_W11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[647%GROUP_COUNT]), .out(W11));
pin_uart #(.NAME("Y1")) pin_Y1_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[648%GROUP_COUNT]), .out(Y1));
pin_uart #(.NAME("Y2")) pin_Y2_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[649%GROUP_COUNT]), .out(Y2));
pin_uart #(.NAME("Y4")) pin_Y4_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[650%GROUP_COUNT]), .out(Y4));
pin_uart #(.NAME("Y6")) pin_Y6_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[651%GROUP_COUNT]), .out(Y6));
pin_uart #(.NAME("Y7")) pin_Y7_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[652%GROUP_COUNT]), .out(Y7));
pin_uart #(.NAME("Y8")) pin_Y8_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[653%GROUP_COUNT]), .out(Y8));
pin_uart #(.NAME("Y9")) pin_Y9_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[654%GROUP_COUNT]), .out(Y9));
pin_uart #(.NAME("Y11")) pin_Y11_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[655%GROUP_COUNT]), .out(Y11));
pin_uart #(.NAME("Y12")) pin_Y12_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[656%GROUP_COUNT]), .out(Y12));
pin_uart #(.NAME("Y13")) pin_Y13_uart_inst (.clk(clk_int), .rst(shift_rst_reg), .shift(shift_reg[657%GROUP_COUNT]), .out(Y13));
endmodule

`resetall
